module MIPS(
    //Input 
    clk,
    rst_n,
    in_valid,
    instruction,
	output_reg,
    //OUTPUT
    out_valid,
    out_1,
	out_2,
	out_3,
	out_4,
	instruction_fail
);

//Input 
input clk;
input rst_n;
input in_valid;
input [31:0] instruction;
input [19:0] output_reg;
//OUTPUT
output logic out_valid, instruction_fail;
output logic [15:0] out_1, out_2, out_3, out_4;

logic [19:0]out,out_reg;
logic[15:0] address[0:5];
logic[15:0] address_reg[0:5];

logic [15:0]in_reg,in;
typedef enum logic [2:0] {IDLE , OUTPUT ,FAIL,WAIT,WAITFAIL,GCD } state;
state curr,next;

logic [15:0]gcda,gcda_reg, gcdb,gcdb_reg;
logic [2:0]Rs , Rt ,Rd; 

logic [2:0]Rd_reg;
logic [15:0]ans,ans_reg;
logic [3:0]shifta,shiftb ,shiftab;
logic in_valid1;
logic a;
always_ff @( posedge clk , negedge rst_n ) begin : state_DFF
    if(!rst_n)begin 
        curr<=IDLE;
    end
    else begin
        curr<=next;
    end
end

always_ff @( posedge clk , negedge rst_n ) begin : address_DFF
    if(!rst_n)begin
        address_reg[0]<=0;
        address_reg[1]<=0;
        address_reg[2]<=0;
        address_reg[3]<=0;
        address_reg[4]<=0;
        address_reg[5]<=0;
        //out_reg<=0;
        //Rd_reg<=0;
        //ans_reg<=0;
    end
    else begin
        address_reg<=address;
        
    end
end

always_comb begin : find_gcd_1
    case (gcda_reg)
        2:a=1;3:a=1;5:a=1;7:a=1;11:a=1;13:a=1;17:a=1;19:a=1;23:a=1;29:a=1;
        31:a=1;37:a=1;41:a=1;43:a=1;47:a=1;53:a=1;59:a=1;61:a=1;67:a=1;71:a=1;
        73:a=1;79:a=1;83:a=1;89:a=1;97:a=1;101:a=1;103:a=1;107:a=1;109:a=1;113:a=1;
        127:a=1;131:a=1;137:a=1;139:a=1;149:a=1;151:a=1;157:a=1;163:a=1;167:a=1;173:a=1;
        179:a=1;181:a=1;191:a=1;193:a=1;197:a=1;199:a=1;211:a=1;223:a=1;227:a=1;229:a=1;
        233:a=1;239:a=1;241:a=1;251:a=1;257:a=1;263:a=1;269:a=1;271:a=1;277:a=1;281:a=1;
        283:a=1;293:a=1;307:a=1;311:a=1;313:a=1;317:a=1;331:a=1;337:a=1;347:a=1;349:a=1;
        353:a=1;359:a=1;367:a=1;373:a=1;379:a=1;383:a=1;389:a=1;397:a=1;401:a=1;409:a=1;
        419:a=1;421:a=1;431:a=1;433:a=1;439:a=1;443:a=1;449:a=1;457:a=1;461:a=1;463:a=1;
        467:a=1;479:a=1;487:a=1;491:a=1;499:a=1;503:a=1;509:a=1;521:a=1;523:a=1;541:a=1;
        547:a=1;557:a=1;563:a=1;569:a=1;571:a=1;577:a=1;587:a=1;593:a=1;599:a=1;601:a=1;
        607:a=1;613:a=1;617:a=1;619:a=1;631:a=1;641:a=1;643:a=1;647:a=1;653:a=1;659:a=1;
        661:a=1;673:a=1;677:a=1;683:a=1;691:a=1;701:a=1;709:a=1;719:a=1;727:a=1;733:a=1;
        739:a=1;743:a=1;751:a=1;757:a=1;761:a=1;769:a=1;773:a=1;787:a=1;797:a=1;809:a=1;
        811:a=1;821:a=1;823:a=1;827:a=1;829:a=1;839:a=1;853:a=1;857:a=1;859:a=1;863:a=1;
        877:a=1;881:a=1;883:a=1;887:a=1;907:a=1;911:a=1;919:a=1;929:a=1;937:a=1;941:a=1;
        947:a=1;953:a=1;967:a=1;971:a=1;977:a=1;983:a=1;991:a=1;997:a=1;1009:a=1;1013:a=1;
        1019:a=1;1021:a=1;1031:a=1;1033:a=1;1039:a=1;1049:a=1;1051:a=1;1061:a=1;1063:a=1;1069:a=1;
        1087:a=1;1091:a=1;1093:a=1;1097:a=1;1103:a=1;1109:a=1;1117:a=1;1123:a=1;1129:a=1;1151:a=1;
        1153:a=1;1163:a=1;1171:a=1;1181:a=1;1187:a=1;1193:a=1;1201:a=1;1213:a=1;1217:a=1;1223:a=1;
        1229:a=1;1231:a=1;1237:a=1;1249:a=1;1259:a=1;1277:a=1;1279:a=1;1283:a=1;1289:a=1;1291:a=1;
        1297:a=1;1301:a=1;1303:a=1;1307:a=1;1319:a=1;1321:a=1;1327:a=1;1361:a=1;1367:a=1;1373:a=1;
        1381:a=1;1399:a=1;1409:a=1;1423:a=1;1427:a=1;1429:a=1;1433:a=1;1439:a=1;1447:a=1;1451:a=1;
        1453:a=1;1459:a=1;1471:a=1;1481:a=1;1483:a=1;1487:a=1;1489:a=1;1493:a=1;1499:a=1;1511:a=1;
        1523:a=1;1531:a=1;1543:a=1;1549:a=1;1553:a=1;1559:a=1;1567:a=1;1571:a=1;1579:a=1;1583:a=1;
        1597:a=1;1601:a=1;1607:a=1;1609:a=1;1613:a=1;1619:a=1;1621:a=1;1627:a=1;1637:a=1;1657:a=1;
        1663:a=1;1667:a=1;1669:a=1;1693:a=1;1697:a=1;1699:a=1;1709:a=1;1721:a=1;1723:a=1;1733:a=1;
        1741:a=1;1747:a=1;1753:a=1;1759:a=1;1777:a=1;1783:a=1;1787:a=1;1789:a=1;1801:a=1;1811:a=1;
        1823:a=1;1831:a=1;1847:a=1;1861:a=1;1867:a=1;1871:a=1;1873:a=1;1877:a=1;1879:a=1;1889:a=1;
        1901:a=1;1907:a=1;1913:a=1;1931:a=1;1933:a=1;1949:a=1;1951:a=1;1973:a=1;1979:a=1;1987:a=1;
        1993:a=1;1997:a=1;1999:a=1;2003:a=1;2011:a=1;2017:a=1;2027:a=1;2029:a=1;2039:a=1;2053:a=1;
        2063:a=1;2069:a=1;2081:a=1;2083:a=1;2087:a=1;2089:a=1;2099:a=1;2111:a=1;2113:a=1;2129:a=1;
        2131:a=1;2137:a=1;2141:a=1;2143:a=1;2153:a=1;2161:a=1;2179:a=1;2203:a=1;2207:a=1;2213:a=1;
        2221:a=1;2237:a=1;2239:a=1;2243:a=1;2251:a=1;2267:a=1;2269:a=1;2273:a=1;2281:a=1;2287:a=1;
        2293:a=1;2297:a=1;2309:a=1;2311:a=1;2333:a=1;2339:a=1;2341:a=1;2347:a=1;2351:a=1;2357:a=1;
        2371:a=1;2377:a=1;2381:a=1;2383:a=1;2389:a=1;2393:a=1;2399:a=1;2411:a=1;2417:a=1;2423:a=1;
        2437:a=1;2441:a=1;2447:a=1;2459:a=1;2467:a=1;2473:a=1;2477:a=1;2503:a=1;2521:a=1;2531:a=1;
        2539:a=1;2543:a=1;2549:a=1;2551:a=1;2557:a=1;2579:a=1;2591:a=1;2593:a=1;2609:a=1;2617:a=1;
        2621:a=1;2633:a=1;2647:a=1;2657:a=1;2659:a=1;2663:a=1;2671:a=1;2677:a=1;2683:a=1;2687:a=1;
        2689:a=1;2693:a=1;2699:a=1;2707:a=1;2711:a=1;2713:a=1;2719:a=1;2729:a=1;2731:a=1;2741:a=1;
        2749:a=1;2753:a=1;2767:a=1;2777:a=1;2789:a=1;2791:a=1;2797:a=1;2801:a=1;2803:a=1;2819:a=1;
        2833:a=1;2837:a=1;2843:a=1;2851:a=1;2857:a=1;2861:a=1;2879:a=1;2887:a=1;2897:a=1;2903:a=1;
        2909:a=1;2917:a=1;2927:a=1;2939:a=1;2953:a=1;2957:a=1;2963:a=1;2969:a=1;2971:a=1;2999:a=1;
        3001:a=1;3011:a=1;3019:a=1;3023:a=1;3037:a=1;3041:a=1;3049:a=1;3061:a=1;3067:a=1;3079:a=1;
        3083:a=1;3089:a=1;3109:a=1;3119:a=1;3121:a=1;3137:a=1;3163:a=1;3167:a=1;3169:a=1;3181:a=1;
        3187:a=1;3191:a=1;3203:a=1;3209:a=1;3217:a=1;3221:a=1;3229:a=1;3251:a=1;3253:a=1;3257:a=1;
        3259:a=1;3271:a=1;3299:a=1;3301:a=1;3307:a=1;3313:a=1;3319:a=1;3323:a=1;3329:a=1;3331:a=1;
        3343:a=1;3347:a=1;3359:a=1;3361:a=1;3371:a=1;3373:a=1;3389:a=1;3391:a=1;3407:a=1;3413:a=1;
        3433:a=1;3449:a=1;3457:a=1;3461:a=1;3463:a=1;3467:a=1;3469:a=1;3491:a=1;3499:a=1;3511:a=1;
        3517:a=1;3527:a=1;3529:a=1;3533:a=1;3539:a=1;3541:a=1;3547:a=1;3557:a=1;3559:a=1;3571:a=1;
        3581:a=1;3583:a=1;3593:a=1;3607:a=1;3613:a=1;3617:a=1;3623:a=1;3631:a=1;3637:a=1;3643:a=1;
        3659:a=1;3671:a=1;3673:a=1;3677:a=1;3691:a=1;3697:a=1;3701:a=1;3709:a=1;3719:a=1;3727:a=1;
        3733:a=1;3739:a=1;3761:a=1;3767:a=1;3769:a=1;3779:a=1;3793:a=1;3797:a=1;3803:a=1;3821:a=1;
        3823:a=1;3833:a=1;3847:a=1;3851:a=1;3853:a=1;3863:a=1;3877:a=1;3881:a=1;3889:a=1;3907:a=1;
        3911:a=1;3917:a=1;3919:a=1;3923:a=1;3929:a=1;3931:a=1;3943:a=1;3947:a=1;3967:a=1;3989:a=1;
        4001:a=1;4003:a=1;4007:a=1;4013:a=1;4019:a=1;4021:a=1;4027:a=1;4049:a=1;4051:a=1;4057:a=1;
        4073:a=1;4079:a=1;4091:a=1;4093:a=1;4099:a=1;4111:a=1;4127:a=1;4129:a=1;4133:a=1;4139:a=1;
        4153:a=1;4157:a=1;4159:a=1;4177:a=1;4201:a=1;4211:a=1;4217:a=1;4219:a=1;4229:a=1;4231:a=1;
        4241:a=1;4243:a=1;4253:a=1;4259:a=1;4261:a=1;4271:a=1;4273:a=1;4283:a=1;4289:a=1;4297:a=1;
        4327:a=1;4337:a=1;4339:a=1;4349:a=1;4357:a=1;4363:a=1;4373:a=1;4391:a=1;4397:a=1;4409:a=1;
        4421:a=1;4423:a=1;4441:a=1;4447:a=1;4451:a=1;4457:a=1;4463:a=1;4481:a=1;4483:a=1;4493:a=1;
        4507:a=1;4513:a=1;4517:a=1;4519:a=1;4523:a=1;4547:a=1;4549:a=1;4561:a=1;4567:a=1;4583:a=1;
        4591:a=1;4597:a=1;4603:a=1;4621:a=1;4637:a=1;4639:a=1;4643:a=1;4649:a=1;4651:a=1;4657:a=1;
        4663:a=1;4673:a=1;4679:a=1;4691:a=1;4703:a=1;4721:a=1;4723:a=1;4729:a=1;4733:a=1;4751:a=1;
        4759:a=1;4783:a=1;4787:a=1;4789:a=1;4793:a=1;4799:a=1;4801:a=1;4813:a=1;4817:a=1;4831:a=1;
        4861:a=1;4871:a=1;4877:a=1;4889:a=1;4903:a=1;4909:a=1;4919:a=1;4931:a=1;4933:a=1;4937:a=1;
        4943:a=1;4951:a=1;4957:a=1;4967:a=1;4969:a=1;4973:a=1;4987:a=1;4993:a=1;4999:a=1;5003:a=1;
        5009:a=1;5011:a=1;5021:a=1;5023:a=1;5039:a=1;5051:a=1;5059:a=1;5077:a=1;5081:a=1;5087:a=1;
        5099:a=1;5101:a=1;5107:a=1;5113:a=1;5119:a=1;5147:a=1;5153:a=1;5167:a=1;5171:a=1;5179:a=1;
        5189:a=1;5197:a=1;5209:a=1;5227:a=1;5231:a=1;5233:a=1;5237:a=1;5261:a=1;5273:a=1;5279:a=1;
        5281:a=1;5297:a=1;5303:a=1;5309:a=1;5323:a=1;5333:a=1;5347:a=1;5351:a=1;5381:a=1;5387:a=1;
        5393:a=1;5399:a=1;5407:a=1;5413:a=1;5417:a=1;5419:a=1;5431:a=1;5437:a=1;5441:a=1;5443:a=1;
        5449:a=1;5471:a=1;5477:a=1;5479:a=1;5483:a=1;5501:a=1;5503:a=1;5507:a=1;5519:a=1;5521:a=1;
        5527:a=1;5531:a=1;5557:a=1;5563:a=1;5569:a=1;5573:a=1;5581:a=1;5591:a=1;5623:a=1;5639:a=1;
        5641:a=1;5647:a=1;5651:a=1;5653:a=1;5657:a=1;5659:a=1;5669:a=1;5683:a=1;5689:a=1;5693:a=1;
        5701:a=1;5711:a=1;5717:a=1;5737:a=1;5741:a=1;5743:a=1;5749:a=1;5779:a=1;5783:a=1;5791:a=1;
        5801:a=1;5807:a=1;5813:a=1;5821:a=1;5827:a=1;5839:a=1;5843:a=1;5849:a=1;5851:a=1;5857:a=1;
        5861:a=1;5867:a=1;5869:a=1;5879:a=1;5881:a=1;5897:a=1;5903:a=1;5923:a=1;5927:a=1;5939:a=1;
        5953:a=1;5981:a=1;5987:a=1;6007:a=1;6011:a=1;6029:a=1;6037:a=1;6043:a=1;6047:a=1;6053:a=1;
        6067:a=1;6073:a=1;6079:a=1;6089:a=1;6091:a=1;6101:a=1;6113:a=1;6121:a=1;6131:a=1;6133:a=1;
        6143:a=1;6151:a=1;6163:a=1;6173:a=1;6197:a=1;6199:a=1;6203:a=1;6211:a=1;6217:a=1;6221:a=1;
        6229:a=1;6247:a=1;6257:a=1;6263:a=1;6269:a=1;6271:a=1;6277:a=1;6287:a=1;6299:a=1;6301:a=1;
        6311:a=1;6317:a=1;6323:a=1;6329:a=1;6337:a=1;6343:a=1;6353:a=1;6359:a=1;6361:a=1;6367:a=1;
        6373:a=1;6379:a=1;6389:a=1;6397:a=1;6421:a=1;6427:a=1;6449:a=1;6451:a=1;6469:a=1;6473:a=1;
        6481:a=1;6491:a=1;6521:a=1;6529:a=1;6547:a=1;6551:a=1;6553:a=1;6563:a=1;6569:a=1;6571:a=1;
        6577:a=1;6581:a=1;6599:a=1;6607:a=1;6619:a=1;6637:a=1;6653:a=1;6659:a=1;6661:a=1;6673:a=1;
        6679:a=1;6689:a=1;6691:a=1;6701:a=1;6703:a=1;6709:a=1;6719:a=1;6733:a=1;6737:a=1;6761:a=1;
        6763:a=1;6779:a=1;6781:a=1;6791:a=1;6793:a=1;6803:a=1;6823:a=1;6827:a=1;6829:a=1;6833:a=1;
        6841:a=1;6857:a=1;6863:a=1;6869:a=1;6871:a=1;6883:a=1;6899:a=1;6907:a=1;6911:a=1;6917:a=1;
        6947:a=1;6949:a=1;6959:a=1;6961:a=1;6967:a=1;6971:a=1;6977:a=1;6983:a=1;6991:a=1;6997:a=1;
        7001:a=1;7013:a=1;7019:a=1;7027:a=1;7039:a=1;7043:a=1;7057:a=1;7069:a=1;7079:a=1;7103:a=1;
        7109:a=1;7121:a=1;7127:a=1;7129:a=1;7151:a=1;7159:a=1;7177:a=1;7187:a=1;7193:a=1;7207:a=1;
        7211:a=1;7213:a=1;7219:a=1;7229:a=1;7237:a=1;7243:a=1;7247:a=1;7253:a=1;7283:a=1;7297:a=1;
        7307:a=1;7309:a=1;7321:a=1;7331:a=1;7333:a=1;7349:a=1;7351:a=1;7369:a=1;7393:a=1;7411:a=1;
        7417:a=1;7433:a=1;7451:a=1;7457:a=1;7459:a=1;7477:a=1;7481:a=1;7487:a=1;7489:a=1;7499:a=1;
        7507:a=1;7517:a=1;7523:a=1;7529:a=1;7537:a=1;7541:a=1;7547:a=1;7549:a=1;7559:a=1;7561:a=1;
        7573:a=1;7577:a=1;7583:a=1;7589:a=1;7591:a=1;7603:a=1;7607:a=1;7621:a=1;7639:a=1;7643:a=1;
        7649:a=1;7669:a=1;7673:a=1;7681:a=1;7687:a=1;7691:a=1;7699:a=1;7703:a=1;7717:a=1;7723:a=1;
        7727:a=1;7741:a=1;7753:a=1;7757:a=1;7759:a=1;7789:a=1;7793:a=1;7817:a=1;7823:a=1;7829:a=1;
        7841:a=1;7853:a=1;7867:a=1;7873:a=1;7877:a=1;7879:a=1;7883:a=1;7901:a=1;7907:a=1;7919:a=1;
        7927:a=1;7933:a=1;7937:a=1;7949:a=1;7951:a=1;7963:a=1;7993:a=1;8009:a=1;8011:a=1;8017:a=1;
        8039:a=1;8053:a=1;8059:a=1;8069:a=1;8081:a=1;8087:a=1;8089:a=1;8093:a=1;8101:a=1;8111:a=1;
        8117:a=1;8123:a=1;8147:a=1;8161:a=1;8167:a=1;8171:a=1;8179:a=1;8191:a=1;8209:a=1;8219:a=1;
        8221:a=1;8231:a=1;8233:a=1;8237:a=1;8243:a=1;8263:a=1;8269:a=1;8273:a=1;8287:a=1;8291:a=1;
        8293:a=1;8297:a=1;8311:a=1;8317:a=1;8329:a=1;8353:a=1;8363:a=1;8369:a=1;8377:a=1;8387:a=1;
        8389:a=1;8419:a=1;8423:a=1;8429:a=1;8431:a=1;8443:a=1;8447:a=1;8461:a=1;8467:a=1;8501:a=1;
        8513:a=1;8521:a=1;8527:a=1;8537:a=1;8539:a=1;8543:a=1;8563:a=1;8573:a=1;8581:a=1;8597:a=1;
        8599:a=1;8609:a=1;8623:a=1;8627:a=1;8629:a=1;8641:a=1;8647:a=1;8663:a=1;8669:a=1;8677:a=1;
        8681:a=1;8689:a=1;8693:a=1;8699:a=1;8707:a=1;8713:a=1;8719:a=1;8731:a=1;8737:a=1;8741:a=1;
        8747:a=1;8753:a=1;8761:a=1;8779:a=1;8783:a=1;8803:a=1;8807:a=1;8819:a=1;8821:a=1;8831:a=1;
        8837:a=1;8839:a=1;8849:a=1;8861:a=1;8863:a=1;8867:a=1;8887:a=1;8893:a=1;8923:a=1;8929:a=1;
        8933:a=1;8941:a=1;8951:a=1;8963:a=1;8969:a=1;8971:a=1;8999:a=1;9001:a=1;9007:a=1;9011:a=1;
        9013:a=1;9029:a=1;9041:a=1;9043:a=1;9049:a=1;9059:a=1;9067:a=1;9091:a=1;9103:a=1;9109:a=1;
        9127:a=1;9133:a=1;9137:a=1;9151:a=1;9157:a=1;9161:a=1;9173:a=1;9181:a=1;9187:a=1;9199:a=1;
        9203:a=1;9209:a=1;9221:a=1;9227:a=1;9239:a=1;9241:a=1;9257:a=1;9277:a=1;9281:a=1;9283:a=1;
        9293:a=1;9311:a=1;9319:a=1;9323:a=1;9337:a=1;9341:a=1;9343:a=1;9349:a=1;9371:a=1;9377:a=1;
        9391:a=1;9397:a=1;9403:a=1;9413:a=1;9419:a=1;9421:a=1;9431:a=1;9433:a=1;9437:a=1;9439:a=1;
        9461:a=1;9463:a=1;9467:a=1;9473:a=1;9479:a=1;9491:a=1;9497:a=1;9511:a=1;9521:a=1;9533:a=1;
        9539:a=1;9547:a=1;9551:a=1;9587:a=1;9601:a=1;9613:a=1;9619:a=1;9623:a=1;9629:a=1;9631:a=1;
        9643:a=1;9649:a=1;9661:a=1;9677:a=1;9679:a=1;9689:a=1;9697:a=1;9719:a=1;9721:a=1;9733:a=1;
        9739:a=1;9743:a=1;9749:a=1;9767:a=1;9769:a=1;9781:a=1;9787:a=1;9791:a=1;9803:a=1;9811:a=1;
        9817:a=1;9829:a=1;9833:a=1;9839:a=1;9851:a=1;9857:a=1;9859:a=1;9871:a=1;9883:a=1;9887:a=1;
        9901:a=1;9907:a=1;9923:a=1;9929:a=1;9931:a=1;9941:a=1;9949:a=1;9967:a=1;9973:a=1;10007:a=1;
        default: a=0;
    endcase
   
end
always_ff @( posedge clk ) begin : gcd_DFF
    gcda_reg<=gcda;
    gcdb_reg<=gcdb;
    out_reg<=out;
    Rd_reg<=Rd;
    ans_reg<=ans;
    in_valid1<=in_valid;
end

always_comb begin : FSM
    
    gcda=0;
    gcdb=0;
    
    Rs=0;
    Rt=0;
    
    shifta=0;
    shifta=0;
    shiftab=0;
    case (curr)
        IDLE:begin
            ans=1;
            address=address_reg;
            out_1=0;
            out_2=0;
            out_3=0;
            out_4=0;
            out_valid=0;
            instruction_fail=0;
            if(in_valid)begin
                out=output_reg;

                case(instruction[25:21])
                    5'b10001:Rs=0;
                    5'b10010:Rs=1;
                    5'b01000:Rs=2;
                    5'b10111:Rs=3;
                    5'b11111:Rs=4;
                    5'b10000:Rs=5;
                    default: Rs=6;
                endcase

                case(instruction[20:16])
                    5'b10001:Rt=0;
                    5'b10010:Rt=1;
                    5'b01000:Rt=2;
                    5'b10111:Rt=3;
                    5'b11111:Rt=4;
                    5'b10000:Rt=5;
                    default: Rt=6;
                endcase

                 case(instruction[15:11])
                    5'b10001:Rd=0;
                    5'b10010:Rd=1;
                    5'b01000:Rd=2;
                    5'b10111:Rd=3;
                    5'b11111:Rd=4;
                    5'b10000:Rd=5;
                    default: Rd=6;
                endcase
                if(instruction[31:26]==6'b000000)begin
                    if(Rt==6||Rs==6||Rd==6)begin
                        next=WAITFAIL;
                    end
                    else begin
                        next=WAIT;
                        case (instruction[6:0])
                            7'b0100000:address[Rd]=(address_reg[Rs])+(address_reg[Rt]);
                            7'b0100100:address[Rd]=(address_reg[Rs])&(address_reg[Rt]);
                            7'b0100101:address[Rd]=(address_reg[Rs])|(address_reg[Rt]);
                            7'b0100111:address[Rd]=~((address_reg[Rs])|(address_reg[Rt]));
                            7'b0000000:address[Rd]=(address_reg[Rt])<<(instruction[10:7]);
                            7'b0000010:address[Rd]=(address_reg[Rt])>>(instruction[10:7]);
                            7'b1111000:begin
                                if(!(address_reg[Rs]&&address_reg[Rt])) next=WAITFAIL;
                                else begin
                                    next=GCD;
                                    if(address_reg[Rs]>address_reg[Rt])begin
                                            gcda=address_reg[Rs];
                                            gcdb=address_reg[Rt];
                                        
                                    end
                                    else begin
                                            gcda=address_reg[Rt];
                                            gcdb=address_reg[Rs];
                                        
                                    end
                                    
                                end
                            end
                            default:next=WAITFAIL; 
                        endcase
                    end
                end
                else if(instruction[31:26]==6'b001000)begin
                    if(Rs==6||Rt==6)begin
                        next=WAITFAIL;
                    end
                    else begin
                        next=WAIT;
                        address[Rt]=address_reg[Rs]+instruction[15:0];
                    end
                end
                else begin
                    next=WAITFAIL;
                end

                
            end
            else begin
                next=IDLE;
                out=0;
                Rd=0;
            end
        end
        
        GCD:begin
            
            out=out_reg;
            out_valid=0;
            instruction_fail=0;
            out_1=0;
            out_2=0;
            out_3=0;
            out_4=0;
            
            address=address_reg;

            

            if(gcdb_reg<=1 || gcdb_reg==gcda_reg || (a&&gcdb_reg!=gcda_reg))begin
                Rd=0;
                ans=0;
                address[Rd_reg]=(gcdb_reg==1 || (a&&gcdb_reg!=gcda_reg))?ans_reg:ans_reg*gcda_reg;
                if(in_valid1)begin
                    next=OUTPUT;
                    out_valid=0;
                    instruction_fail=0;
                    out_1=0;
                    out_2=0;
                    out_3=0;
                    out_4=0;
                end
                else begin
                    
                    next=IDLE;              
                    out_valid=1;
                    instruction_fail=0;
                    case(out_reg[19:15])
                        5'b10001:out_4=address[0];
                        5'b10010:out_4=address[1];
                        5'b01000:out_4=address[2];
                        5'b10111:out_4=address[3];
                        5'b11111:out_4=address[4];
                        5'b10000:out_4=address[5];
                        default: out_4=0;
                    endcase

                    case(out_reg[14:10])
                        5'b10001:out_3=address[0];
                        5'b10010:out_3=address[1];
                        5'b01000:out_3=address[2];
                        5'b10111:out_3=address[3];
                        5'b11111:out_3=address[4];
                        5'b10000:out_3=address[5];
                        default: out_3=0;
                    endcase

                    case(out_reg[9:5])
                        5'b10001:out_2=address[0];
                        5'b10010:out_2=address[1];
                        5'b01000:out_2=address[2];
                        5'b10111:out_2=address[3];
                        5'b11111:out_2=address[4];
                        5'b10000:out_2=address[5];
                        default: out_2=0;
                    endcase

                    case(out_reg[4:0])
                        5'b10001:out_1=address[0];
                        5'b10010:out_1=address[1];
                        5'b01000:out_1=address[2];
                        5'b10111:out_1=address[3];
                        5'b11111:out_1=address[4];
                        5'b10000:out_1=address[5];
                        default: out_1=0;
                    endcase      
                    
                end

            end
            else if(gcda_reg[0]==0||gcdb_reg[0]==0)begin
                next=GCD;
                Rd=Rd_reg;
                casez (gcda_reg)
                    16'b??????????????10:shifta= 1;
                    16'b?????????????100:shifta= 2;
                    16'b????????????1000:shifta= 3;
                    16'b???????????10000:shifta= 4;
                    16'b??????????100000:shifta= 5;
                    16'b?????????1000000:shifta= 6;
                    16'b????????10000000:shifta= 7;
                    16'b???????100000000:shifta= 8;
                    16'b??????1000000000:shifta=9; 
                    16'b?????10000000000:shifta=10; 
                    16'b????100000000000:shifta=11; 
                    16'b???1000000000000:shifta=12; 
                    16'b??10000000000000:shifta=13; 
                    16'b?100000000000000:shifta=14; 
                    16'b1000000000000000:shifta=15; 
                    default: shifta=0;
                endcase
                casez (gcdb_reg)
                    16'b??????????????10:shiftb= 1; 
                    16'b?????????????100:shiftb= 2;  
                    16'b????????????1000:shiftb= 3;  
                    16'b???????????10000:shiftb= 4;  
                    16'b??????????100000:shiftb= 5;  
                    16'b?????????1000000:shiftb= 6;  
                    16'b????????10000000:shiftb= 7;  
                    16'b???????100000000:shiftb= 8;  
                    16'b??????1000000000:shiftb=9;   
                    16'b?????10000000000:shiftb=10; 
                    16'b????100000000000:shiftb=11;
                    16'b???1000000000000:shiftb=12;
                    16'b??10000000000000:shiftb=13;
                    16'b?100000000000000:shiftb=14;
                    16'b1000000000000000:shiftb=15;
                    default: shiftb=0;
                endcase
                ans=(shifta<shiftb)?(ans_reg<<shifta):(ans_reg<<shiftb);
                if(gcda_reg>>shifta > gcdb_reg>>shiftb)begin
                    gcda=gcda_reg>>shifta;
                    gcdb=gcdb_reg>>shiftb;
                end
                else begin
                    gcdb=gcda_reg>>shifta;
                    gcda=gcdb_reg>>shiftb;
                end
            end
                
        
           
            
            else begin
                next=GCD;
                Rd=Rd_reg;
                ans=ans_reg;
                casez (gcda_reg-gcdb_reg)
                    16'b??????????????10:shiftab= 1; 
                    16'b?????????????100:shiftab= 2;  
                    16'b????????????1000:shiftab= 3;  
                    16'b???????????10000:shiftab= 4;  
                    16'b??????????100000:shiftab= 5;  
                    16'b?????????1000000:shiftab= 6;  
                    16'b????????10000000:shiftab= 7;  
                    16'b???????100000000:shiftab= 8;  
                    16'b??????1000000000:shiftab=9;   
                    16'b?????10000000000:shiftab=10; 
                    16'b????100000000000:shiftab=11;
                    16'b???1000000000000:shiftab=12;
                    16'b??10000000000000:shiftab=13;
                    16'b?100000000000000:shiftab=14;
                    16'b1000000000000000:shiftab=15;
                    default: shiftab=0;
                endcase
                if((gcda_reg-gcdb_reg)>>shiftab>=gcdb_reg)begin
                    gcda=(gcda_reg-gcdb_reg)>>shiftab;
                    gcdb=gcdb_reg;
                end
                else begin
                    gcdb=(gcda_reg-gcdb_reg)>>shiftab;
                    gcda=gcdb_reg;
                end     
            end       
        
        end
        WAIT:begin
             Rd=0;
            ans=1;
            instruction_fail=0;
            out_valid=0;
            out=out_reg;
            out_1=0;
            out_2=0;
            out_3=0;
            out_4=0;
            address=address_reg;
            next=OUTPUT;
        end
        WAITFAIL:begin
             Rd=0;
            ans=1;
            instruction_fail=0;
            out_valid=0;
            out_1=0;
            out_2=0;
            out_3=0;
            out_4=0;
            out=0;
            address=address_reg;
            next=FAIL;
        end
        OUTPUT:begin
             Rd=0;
            ans=1;
            instruction_fail=0;
            out=0;
            address=address_reg;
            out_valid=1;
            case(out_reg[19:15])
                    5'b10001:out_4=address[0];
                    5'b10010:out_4=address[1];
                    5'b01000:out_4=address[2];
                    5'b10111:out_4=address[3];
                    5'b11111:out_4=address[4];
                    5'b10000:out_4=address[5];
                    default: out_4=0;
                endcase

                case(out_reg[14:10])
                    5'b10001:out_3=address[0];
                    5'b10010:out_3=address[1];
                    5'b01000:out_3=address[2];
                    5'b10111:out_3=address[3];
                    5'b11111:out_3=address[4];
                    5'b10000:out_3=address[5];
                    default: out_3=0;
                endcase

                case(out_reg[9:5])
                    5'b10001:out_2=address[0];
                    5'b10010:out_2=address[1];
                    5'b01000:out_2=address[2];
                    5'b10111:out_2=address[3];
                    5'b11111:out_2=address[4];
                    5'b10000:out_2=address[5];
                    default: out_2=0;
                endcase

                case(out_reg[4:0])
                    5'b10001:out_1=address[0];
                    5'b10010:out_1=address[1];
                    5'b01000:out_1=address[2];
                    5'b10111:out_1=address[3];
                    5'b11111:out_1=address[4];
                    5'b10000:out_1=address[5];
                    default: out_1=0;
                endcase      
            next=IDLE;
        end
        FAIL:begin
             Rd=0;
            ans=1;
            out=0;
            out_1=0;
            out_2=0;
            out_3=0;
            out_4=0;
            address=address_reg;
            out_valid=1;
            instruction_fail=1;
            next=IDLE;
        end
        default:begin
            Rd=0;
            ans=1;
            instruction_fail=0;
            out_valid=0;
            out_1=0;
            out_2=0;
            out_3=0;
            out_4=0;
            out=0;
            address=address_reg;
            next=IDLE;
        end
    endcase
end

endmodule